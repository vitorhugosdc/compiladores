Main{
    main(){
        Teste t;
        t.var1=1.0;
        t.var2;
        t.var5;
        t.funcao2();

        
    }
}